// ADC.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module ADC (
		input  wire        clk_clk,                              //                    clk.clk
		output wire        mm_bridge_0_s0_waitrequest,           //         mm_bridge_0_s0.waitrequest
		output wire [15:0] mm_bridge_0_s0_readdata,              //                       .readdata
		output wire        mm_bridge_0_s0_readdatavalid,         //                       .readdatavalid
		input  wire [0:0]  mm_bridge_0_s0_burstcount,            //                       .burstcount
		input  wire [15:0] mm_bridge_0_s0_writedata,             //                       .writedata
		input  wire [9:0]  mm_bridge_0_s0_address,               //                       .address
		input  wire        mm_bridge_0_s0_write,                 //                       .write
		input  wire        mm_bridge_0_s0_read,                  //                       .read
		input  wire [1:0]  mm_bridge_0_s0_byteenable,            //                       .byteenable
		input  wire        mm_bridge_0_s0_debugaccess,           //                       .debugaccess
		output wire        modular_adc_0_response_valid,         // modular_adc_0_response.valid
		output wire [4:0]  modular_adc_0_response_channel,       //                       .channel
		output wire [11:0] modular_adc_0_response_data,          //                       .data
		output wire        modular_adc_0_response_startofpacket, //                       .startofpacket
		output wire        modular_adc_0_response_endofpacket,   //                       .endofpacket
		input  wire        reset_reset_n                         //                  reset.reset_n
	);

	wire         altpll_0_c0_clk;                                         // altpll_0:c0 -> modular_adc_0:adc_pll_clock_clk
	wire         altpll_0_locked_conduit_export;                          // altpll_0:locked -> modular_adc_0:adc_pll_locked_export
	wire         mm_bridge_0_m0_waitrequest;                              // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [15:0] mm_bridge_0_m0_readdata;                                 // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                              // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [9:0] mm_bridge_0_m0_address;                                  // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                     // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire   [1:0] mm_bridge_0_m0_byteenable;                               // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                            // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [15:0] mm_bridge_0_m0_writedata;                                // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                    // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                               // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire  [31:0] master_0_master_readdata;                                // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                             // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                 // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                    // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                              // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                           // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                   // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                               // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_readdata;  // modular_adc_0:sequencer_csr_readdata -> mm_interconnect_0:modular_adc_0_sequencer_csr_readdata
	wire   [0:0] mm_interconnect_0_modular_adc_0_sequencer_csr_address;   // mm_interconnect_0:modular_adc_0_sequencer_csr_address -> modular_adc_0:sequencer_csr_address
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_read;      // mm_interconnect_0:modular_adc_0_sequencer_csr_read -> modular_adc_0:sequencer_csr_read
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_write;     // mm_interconnect_0:modular_adc_0_sequencer_csr_write -> modular_adc_0:sequencer_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_writedata; // mm_interconnect_0:modular_adc_0_sequencer_csr_writedata -> modular_adc_0:sequencer_csr_writedata
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [altpll_0:reset, mm_bridge_0:reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, modular_adc_0:reset_sink_reset_n]

	ADC_altpll_0 altpll_0 (
		.clk                (clk_clk),                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (altpll_0_c0_clk),                //                    c0.clk
		.locked             (altpll_0_locked_conduit_export), //        locked_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.c1                 (),                               //           (terminated)
		.c2                 (),                               //           (terminated)
		.c3                 (),                               //           (terminated)
		.c4                 (),                               //           (terminated)
		.areset             (1'b0),                           //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (3'b000),                         //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	ADC_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (16),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mm_bridge_0_s0_waitrequest),     //    s0.waitrequest
		.s0_readdata      (mm_bridge_0_s0_readdata),        //      .readdata
		.s0_readdatavalid (mm_bridge_0_s0_readdatavalid),   //      .readdatavalid
		.s0_burstcount    (mm_bridge_0_s0_burstcount),      //      .burstcount
		.s0_writedata     (mm_bridge_0_s0_writedata),       //      .writedata
		.s0_address       (mm_bridge_0_s0_address),         //      .address
		.s0_write         (mm_bridge_0_s0_write),           //      .write
		.s0_read          (mm_bridge_0_s0_read),            //      .read
		.s0_byteenable    (mm_bridge_0_s0_byteenable),      //      .byteenable
		.s0_debugaccess   (mm_bridge_0_s0_debugaccess),     //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //      .address
		.m0_write         (mm_bridge_0_m0_write),           //      .write
		.m0_read          (mm_bridge_0_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),     //      .debugaccess
		.s0_response      (),                               // (terminated)
		.m0_response      (2'b00)                           // (terminated)
	);

	ADC_modular_adc_0 #(
		.is_this_first_or_second_adc (1)
	) modular_adc_0 (
		.clock_clk               (clk_clk),                                                 //          clock.clk
		.reset_sink_reset_n      (~rst_controller_reset_out_reset),                         //     reset_sink.reset_n
		.adc_pll_clock_clk       (altpll_0_c0_clk),                                         //  adc_pll_clock.clk
		.adc_pll_locked_export   (altpll_0_locked_conduit_export),                          // adc_pll_locked.export
		.sequencer_csr_address   (mm_interconnect_0_modular_adc_0_sequencer_csr_address),   //  sequencer_csr.address
		.sequencer_csr_read      (mm_interconnect_0_modular_adc_0_sequencer_csr_read),      //               .read
		.sequencer_csr_write     (mm_interconnect_0_modular_adc_0_sequencer_csr_write),     //               .write
		.sequencer_csr_writedata (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata), //               .writedata
		.sequencer_csr_readdata  (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),  //               .readdata
		.response_valid          (modular_adc_0_response_valid),                            //       response.valid
		.response_channel        (modular_adc_0_response_channel),                          //               .channel
		.response_data           (modular_adc_0_response_data),                             //               .data
		.response_startofpacket  (modular_adc_0_response_startofpacket),                    //               .startofpacket
		.response_endofpacket    (modular_adc_0_response_endofpacket)                       //               .endofpacket
	);

	ADC_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                 //                                clk_0_clk.clk
		.master_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                          // master_0_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                          //  mm_bridge_0_reset_reset_bridge_in_reset.reset
		.master_0_master_address                        (master_0_master_address),                                 //                          master_0_master.address
		.master_0_master_waitrequest                    (master_0_master_waitrequest),                             //                                         .waitrequest
		.master_0_master_byteenable                     (master_0_master_byteenable),                              //                                         .byteenable
		.master_0_master_read                           (master_0_master_read),                                    //                                         .read
		.master_0_master_readdata                       (master_0_master_readdata),                                //                                         .readdata
		.master_0_master_readdatavalid                  (master_0_master_readdatavalid),                           //                                         .readdatavalid
		.master_0_master_write                          (master_0_master_write),                                   //                                         .write
		.master_0_master_writedata                      (master_0_master_writedata),                               //                                         .writedata
		.mm_bridge_0_m0_address                         (mm_bridge_0_m0_address),                                  //                           mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                     (mm_bridge_0_m0_waitrequest),                              //                                         .waitrequest
		.mm_bridge_0_m0_burstcount                      (mm_bridge_0_m0_burstcount),                               //                                         .burstcount
		.mm_bridge_0_m0_byteenable                      (mm_bridge_0_m0_byteenable),                               //                                         .byteenable
		.mm_bridge_0_m0_read                            (mm_bridge_0_m0_read),                                     //                                         .read
		.mm_bridge_0_m0_readdata                        (mm_bridge_0_m0_readdata),                                 //                                         .readdata
		.mm_bridge_0_m0_readdatavalid                   (mm_bridge_0_m0_readdatavalid),                            //                                         .readdatavalid
		.mm_bridge_0_m0_write                           (mm_bridge_0_m0_write),                                    //                                         .write
		.mm_bridge_0_m0_writedata                       (mm_bridge_0_m0_writedata),                                //                                         .writedata
		.mm_bridge_0_m0_debugaccess                     (mm_bridge_0_m0_debugaccess),                              //                                         .debugaccess
		.modular_adc_0_sequencer_csr_address            (mm_interconnect_0_modular_adc_0_sequencer_csr_address),   //              modular_adc_0_sequencer_csr.address
		.modular_adc_0_sequencer_csr_write              (mm_interconnect_0_modular_adc_0_sequencer_csr_write),     //                                         .write
		.modular_adc_0_sequencer_csr_read               (mm_interconnect_0_modular_adc_0_sequencer_csr_read),      //                                         .read
		.modular_adc_0_sequencer_csr_readdata           (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),  //                                         .readdata
		.modular_adc_0_sequencer_csr_writedata          (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata)  //                                         .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
